`ifndef ENUM_SVH
`define ENUM_SVH

typedef enum bit[1:0] { ADD, SUB, BITWISE_INVERT, REDUCTION } opcode_e;

`endif